// a testing package for testing tag cache

`include "config.svh"

package cache_pkg;

   // definition of cache blocks
`include "packet.svh"

   // definition of cache
`include "cache.svh"

   // definition of a processor
`include "processor.svh"


endpackage // cache_pkg
   
