// define all macros

`define LNEndpoints  2

`define TLAddrBits 26

`define TLClientXactIdBits 3

`define TLMasterXactIdBits 1;

`define TLDataBits 544

`define acquireTypeWidth 3

`define TLWriteMaskBits 6

`define TLWordAddrBits 3

`define TLAtomicOpBits 4

`define MIFAddrBits

`define MIFTagBits
 
`define MIFDataBits
