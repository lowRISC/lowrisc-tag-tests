// define the packets used by caches

class acquire;

   rand 
